LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY seg IS
PORT (a:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
     led7s: OUT STD_LOGIC_VECTOR( 6 DOWNTO 0));
END seg;
ARCHITECTURE bhv OF seg IS
BEGIN
PROCESS (a)
BEGIN
IF a= "0000" THEN led7s <= NOT"0111111" ; --共阴极, g a
ELSIF a="0001" THEN led7s <= NOT"0000110";
ELSIF a="0010" THEN led7s <= NOT"1011011";
ELSIF a="0011" THEN led7s <= NOT"1001111";
ELSIF a="0100" THEN led7s <= NOT"1100110";
ELSIF a="0101" THEN led7s <= NOT"1101101";
ELSIF a="0110" THEN led7s <= NOT"1111101";
ELSIF a="0111" THEN led7s <= NOT"0000111";
ELSIF a="1000" THEN led7s <= NOT"1111111";
ELSIF a="1001" THEN led7s <= NOT"1101111";
ELSE led7s<="0000000";
END IF;
END PROCESS;
END;